`timescale 1ns/1ns

module InstructionMemory(
    input[31:0] addr,
    output[31:0] inst_out
);
    reg[7:0] mem[0:1023] ;

	wire[9:0] address;
	assign address = addr[9:0];
  	assign inst_out = {mem[address], mem[address + 1], mem[address + 2], mem[address + 3]} ;
	/*
	always @(posedge clk) begin
		inst_out <= {mem[address], mem[address + 1], mem[address + 2], mem[address + 3]} ;
	end*/
	initial begin
		for ( integer i = 0 ; i < 1024 ; i = i + 1) begin
	    	mem[i] = 8'b0 ;
		end
		{mem[ 0], mem[ 0 + 1], mem[ 0 + 2], mem[ 0 + 3]} = { 6'b100011, 5'b00001, 5'b00010, 5'b00000, 5'b00000, 6'b000000 } ; // LW  R2, R1, 0  -> R2 =  5
		{mem[ 4], mem[ 4 + 1], mem[ 4 + 2], mem[ 4 + 3]} = { 6'b100011, 5'b00001, 5'b00011, 5'b00000, 5'b00000, 6'b000001 } ; // LW  R3, R1, 1  -> R3 = 10
		{mem[ 8], mem[ 8 + 1], mem[ 8 + 2], mem[ 8 + 3]} = { 6'b100011, 5'b00001, 5'b00100, 5'b00000, 5'b00000, 6'b000010 } ; // LW  R4, R1, 2  -> R4 = 1
		{mem[12], mem[12 + 1], mem[12 + 2], mem[12 + 3]} = { 6'b100011, 5'b00001, 5'b00101, 5'b00000, 5'b00000, 6'b000011 } ; // LW  R5, R1, 3  -> R5 = 20
		{mem[16], mem[16 + 1], mem[16 + 2], mem[16 + 3]} = { 6'b100011, 5'b00001, 5'b00110, 5'b00000, 5'b00000, 6'b000100 } ; // LW  R6, R1, 4  -> R6 = 25

		{mem[20], mem[20 + 1], mem[20 + 2], mem[20 + 3]} = { 6'b000000, 5'b00010, 5'b00011, 5'b00111, 5'b00000, 6'b100000 } ; // ADD R7, R2, R3 -> R7 = 15
		{mem[24], mem[24 + 1], mem[24 + 2], mem[24 + 3]} = { 6'b000000, 5'b00111, 5'b00100, 5'b00111, 5'b00000, 6'b100000 } ; // ADD R7, R7, R4 -> R7 = 16
		{mem[28], mem[28 + 1], mem[28 + 2], mem[28 + 3]} = { 6'b000000, 5'b00111, 5'b00101, 5'b00111, 5'b00000, 6'b100000 } ; // ADD R7, R7, R5 -> R7 = 36
		{mem[32], mem[32 + 1], mem[32 + 2], mem[32 + 3]} = { 6'b000000, 5'b00111, 5'b00110, 5'b00111, 5'b00000, 6'b100000 } ; // ADD R7, R7, R6 -> R7 = 61
		{mem[36], mem[36 + 1], mem[36 + 2], mem[36 + 3]} = { 6'b000000, 5'b00111, 5'b00110, 5'b01000, 5'b00000, 6'b100000 } ; // ADD R8, R7, R6 -> R8 = 86
		{mem[40], mem[40 + 1], mem[40 + 2], mem[40 + 3]} = { 6'b000000, 5'b00111, 5'b01000, 5'b01001, 5'b00000, 6'b100000 } ; // ADD R9, R7, R8 -> R9 = 147
		{mem[44], mem[44 + 1], mem[44 + 2], mem[44 + 3]} = { 6'b000000, 5'b01001, 5'b01000, 5'b01010, 5'b00000, 6'b100010 } ; // SUB R10, R9, R8 -> R10 = 61

		{mem[48], mem[48 + 1], mem[48 + 2], mem[48 + 3]} = { 6'b100011, 5'b00001, 5'b01011, 5'b00000, 5'b00000, 6'b000100 } ; // LW  R11, R1, 4 -> R11 = 25
		{mem[52], mem[52 + 1], mem[52 + 2], mem[52 + 3]} = { 6'b000000, 5'b01001, 5'b01011, 5'b01100, 5'b00000, 6'b100000 } ; // ADD R12, R9, R11 -> R12 = 172
		{mem[56], mem[56 + 1], mem[56 + 2], mem[56 + 3]} = { 6'b101011, 5'b00001, 5'b01100, 5'b00000, 5'b00000, 6'b010000 } ; // SW  R12, R1, 128 -> MEM[16] = 172
		{mem[60], mem[60 + 1], mem[60 + 2], mem[60 + 3]} = { 6'b000000, 5'b01001, 5'b01011, 5'b01101, 5'b00000, 6'b100000 } ; // ADD R13, R9, R11 -> R13 = 172

		{mem[64], mem[64 + 1], mem[64 + 2], mem[64 + 3]} = { 6'b000000, 5'b01001, 5'b01011, 5'b01110, 5'b00000, 6'b101010 } ; // SLT R14, R9, R11 -> R14 = 0
		{mem[68], mem[68 + 1], mem[68 + 2], mem[68 + 3]} = { 6'b000000, 5'b01011, 5'b01001, 5'b01111, 5'b00000, 6'b101010 } ; // SLT R15, R11, R9 -> R15 = 1

		{mem[72], mem[72 + 1], mem[72 + 2], mem[72 + 3]} = { 6'b000000, 5'b01110, 5'b01001, 5'b10000, 5'b00000, 6'b100101 } ; // OR  R16, R14, R9 -> R16 = R9
		{mem[76], mem[76 + 1], mem[76 + 2], mem[76 + 3]} = { 6'b000000, 5'b01001, 5'b01010, 5'b10001, 5'b00000, 6'b100100 } ; // AND R17, R9, R10 -> R17 = 147 & 61 = 17

		{mem[80], mem[80 + 1], mem[80 + 2], mem[80 + 3]} = { 6'b000010, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 6'b010110 } ; // J 22 -> 88

		{mem[84], mem[84 + 1], mem[84 + 2], mem[84 + 3]} = { 6'b000000, 5'b01011, 5'b01001, 5'b10010, 5'b00000, 6'b101010 } ; // SLT R18, R11, R9 -> R18 != 1 -> jump
		{mem[88], mem[88 + 1], mem[88 + 2], mem[88 + 3]} = { 6'b000000, 5'b01011, 5'b01001, 5'b10011, 5'b00000, 6'b101010 } ; // SLT R19, R11, R9 -> R19 = 1


		{mem[92], mem[92 + 1], mem[92 + 2], mem[92 + 3]} = { 6'b000100, 5'b00001, 5'b00010, 5'b00000, 5'b00000, 6'b000001 } ; // BEQ R1,R2

		{mem[96 ], mem[96  + 1], mem[96 +  2], mem[96 +  3]} = { 6'b000000, 5'b01011, 5'b01001, 5'b10100, 5'b00000, 6'b101010 } ; // SLT R20, R11, R9 -> R20 = 1
		{mem[100], mem[100 + 1], mem[100 + 2], mem[100 + 3]} = { 6'b000000, 5'b01011, 5'b01001, 5'b10101, 5'b00000, 6'b101010 } ; // SLT R21, R11, R9 -> R21 = 1

		{mem[104], mem[104 + 1], mem[104 + 2], mem[104 + 3]} = { 6'b000101, 5'b00001, 5'b00010, 5'b00000, 5'b00000, 6'b000001 } ; // BNE R1,R2

		{mem[108], mem[108 + 1], mem[108 + 2], mem[108 + 3]} = { 6'b000000, 5'b01011, 5'b01001, 5'b10110, 5'b00000, 6'b101010 } ; // SLT R22, R11, R9 -> R22 != 1
		{mem[112], mem[112 + 1], mem[112 + 2], mem[112 + 3]} = { 6'b000000, 5'b01011, 5'b01001, 5'b10111, 5'b00000, 6'b101010 } ; // SLT R23, R11, R9 -> R23 = 1

		{mem[116], mem[116 + 1], mem[116 + 2], mem[116 + 3]} = { 6'b000000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 6'b000000 } ; // NOP
		{mem[120], mem[120 + 1], mem[120 + 2], mem[120 + 3]} = { 6'b000000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 6'b000000 } ; // NOP
		{mem[124], mem[124 + 1], mem[124 + 2], mem[124 + 3]} = { 6'b000000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 6'b000000 } ; // NOP

		{mem[128], mem[128 + 1], mem[128 + 2], mem[128 + 3]} = { 6'b000101, 5'b00001, 5'b10111, 5'b00000, 5'b00000, 6'b000001 } ; // BNE R1,R23

		{mem[132], mem[132 + 1], mem[132 + 2], mem[132 + 3]} = { 6'b000000, 5'b01011, 5'b01001, 5'b11000, 5'b00000, 6'b101010 } ; // SLT R24, R11, R9 -> R24 != 1
		{mem[136], mem[136 + 1], mem[136 + 2], mem[136 + 3]} = { 6'b000000, 5'b01011, 5'b01001, 5'b11001, 5'b00000, 6'b101010 } ; // SLT R25, R11, R9 -> R25 = 1


	end
endmodule
