`timescale 1ns/1ns

module InstructionMemory(
    input[31:0] addr,
    output[31:0] inst_out
);
    reg[7:0] mem[0:1023] ;

	wire[9:0] address;
	assign address = addr[9:0];
  	assign inst_out = {mem[address], mem[address + 1], mem[address + 2], mem[address + 3]} ;
	/*
	always @(posedge clk) begin
		inst_out <= {mem[address], mem[address + 1], mem[address + 2], mem[address + 3]} ;
	end*/
	initial begin
		for ( integer i = 0 ; i < 1024 ; i = i + 1) begin
	    	mem[i] = 8'b0 ;
		end
		{mem[ 0], mem[ 0 + 1], mem[ 0 + 2], mem[ 0 + 3]} = { 6'b100011, 5'b00001, 5'b00010, 5'b00000, 5'b00000, 6'b000000 } ; // LW  R2, R1, 0  -> R2 =  5
		{mem[ 4], mem[ 4 + 1], mem[ 4 + 2], mem[ 4 + 3]} = { 6'b100011, 5'b00001, 5'b00011, 5'b00000, 5'b00000, 6'b000001 } ; // LW  R3, R1, 1  -> R3 = 10
		{mem[ 8], mem[ 8 + 1], mem[ 8 + 2], mem[ 8 + 3]} = { 6'b100011, 5'b00001, 5'b00100, 5'b00000, 5'b00000, 6'b000010 } ; // LW  R4, R1, 2  -> R4 = 15
		{mem[12], mem[12 + 1], mem[12 + 2], mem[12 + 3]} = { 6'b100011, 5'b00001, 5'b00101, 5'b00000, 5'b00000, 6'b000011 } ; // LW  R5, R1, 3  -> R5 = 20
		{mem[16], mem[16 + 1], mem[16 + 2], mem[16 + 3]} = { 6'b100011, 5'b00001, 5'b00110, 5'b00000, 5'b00000, 6'b000100 } ; // LW  R6, R1, 4  -> R6 = 25

		{mem[20], mem[20 + 1], mem[20 + 2], mem[20 + 3]} = { 6'b000000, 5'b00010, 5'b00011, 5'b00111, 5'b00000, 6'b100000 } ; // ADD R7, R2, R3 -> R7 = 15
		{mem[24], mem[24 + 1], mem[24 + 2], mem[24 + 3]} = { 6'b000000, 5'b00111, 5'b00100, 5'b00111, 5'b00000, 6'b100000 } ; // ADD R7, R7, R4 -> R7 = 30
		{mem[28], mem[28 + 1], mem[28 + 2], mem[28 + 3]} = { 6'b000000, 5'b00111, 5'b00101, 5'b00111, 5'b00000, 6'b100000 } ; // ADD R7, R7, R5 -> R7 = 50
		{mem[32], mem[32 + 1], mem[32 + 2], mem[32 + 3]} = { 6'b000000, 5'b00111, 5'b00110, 5'b00111, 5'b00000, 6'b100000 } ; // ADD R7, R7, R6 -> R7 = 75
		{mem[36], mem[36 + 1], mem[36 + 2], mem[36 + 3]} = { 6'b000000, 5'b00111, 5'b00110, 5'b01000, 5'b00000, 6'b100000 } ; // ADD R8, R7, R6 -> R8 = 100
		{mem[40], mem[40 + 1], mem[40 + 2], mem[40 + 3]} = { 6'b000000, 5'b00111, 5'b01000, 5'b01001, 5'b00000, 6'b100000 } ; // ADD R9, R7, R8 -> R9 = 175
		{mem[44], mem[44 + 1], mem[44 + 2], mem[44 + 3]} = { 6'b000000, 5'b01001, 5'b01000, 5'b01010, 5'b00000, 6'b100010 } ; // SUB R10, R9, R8 -> R10 = 75

		{mem[48], mem[48 + 1], mem[48 + 2], mem[48 + 3]} = { 6'b100011, 5'b00001, 5'b01011, 5'b00000, 5'b00000, 6'b000100 } ; // LW  R11, R1, 4 -> R11 = 25
		{mem[52], mem[52 + 1], mem[52 + 2], mem[52 + 3]} = { 6'b000000, 5'b01001, 5'b01011, 5'b01100, 5'b00000, 6'b100000 } ; // ADD R12, R9, R11 -> R12 = 200
	end
endmodule
